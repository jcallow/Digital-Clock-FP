// CPU_Final_Project.v

// Generated using ACDS version 13.1 162 at 2014.06.14.08:55:10

`timescale 1 ps / 1 ps
module CPU_Final_Project (
		input  wire        clk_clk,                           //                        clk.clk
		output wire [12:0] sram_wire_addr,                    //                  sram_wire.addr
		output wire [1:0]  sram_wire_ba,                      //                           .ba
		output wire        sram_wire_cas_n,                   //                           .cas_n
		output wire        sram_wire_cke,                     //                           .cke
		output wire        sram_wire_cs_n,                    //                           .cs_n
		inout  wire [31:0] sram_wire_dq,                      //                           .dq
		output wire [3:0]  sram_wire_dqm,                     //                           .dqm
		output wire        sram_wire_ras_n,                   //                           .ras_n
		output wire        sram_wire_we_n,                    //                           .we_n
		output wire [7:0]  ledg_external_connection_export,   //   ledg_external_connection.export
		output wire [9:0]  ledr_external_connection_export,   //   ledr_external_connection.export
		input  wire [9:0]  switch_external_connection_export, // switch_external_connection.export
		input  wire [3:0]  btn_external_connection_export,    //    btn_external_connection.export
		input  wire        reset_reset_n,                     //                      reset.reset_n
		output wire        lcd_16207_RS,                      //                  lcd_16207.RS
		output wire        lcd_16207_RW,                      //                           .RW
		inout  wire [7:0]  lcd_16207_data,                    //                           .data
		output wire        lcd_16207_E,                       //                           .E
		output wire        sdram_clk_clk,                     //                  sdram_clk.clk
		output wire [14:0] clock_set_ext_export,              //              clock_set_ext.export
		input  wire [13:0] clock_get_ext_export               //              clock_get_ext.export
	);

	wire         clocks_sys_clk_clk;                                        // clocks:sys_clk -> [btn:clk, clock_get:clk, clock_set:clk, cpu:clk, irq_mapper:clk, jtag_uart:clk, lcd_16207_0:clk, ledg:clk, ledr:clk, mm_interconnect_0:clocks_sys_clk_clk, rst_controller:clk, sram:clk, switch:clk, sysid:clock, timer_0:clk]
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [27:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                               // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                       // mm_interconnect_0:ledg_s1_writedata -> ledg:writedata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                         // mm_interconnect_0:ledg_s1_address -> ledg:address
	wire         mm_interconnect_0_ledg_s1_chipselect;                      // mm_interconnect_0:ledg_s1_chipselect -> ledg:chipselect
	wire         mm_interconnect_0_ledg_s1_write;                           // mm_interconnect_0:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                        // ledg:readdata -> mm_interconnect_0:ledg_s1_readdata
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                       // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                         // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_chipselect;                      // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire         mm_interconnect_0_ledr_s1_write;                           // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                        // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                    // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                      // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                   // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                        // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                     // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire  [31:0] mm_interconnect_0_clock_set_s1_writedata;                  // mm_interconnect_0:clock_set_s1_writedata -> clock_set:writedata
	wire   [1:0] mm_interconnect_0_clock_set_s1_address;                    // mm_interconnect_0:clock_set_s1_address -> clock_set:address
	wire         mm_interconnect_0_clock_set_s1_chipselect;                 // mm_interconnect_0:clock_set_s1_chipselect -> clock_set:chipselect
	wire         mm_interconnect_0_clock_set_s1_write;                      // mm_interconnect_0:clock_set_s1_write -> clock_set:write_n
	wire  [31:0] mm_interconnect_0_clock_set_s1_readdata;                   // clock_set:readdata -> mm_interconnect_0:clock_set_s1_readdata
	wire   [1:0] mm_interconnect_0_clock_get_s1_address;                    // mm_interconnect_0:clock_get_s1_address -> clock_get:address
	wire  [31:0] mm_interconnect_0_clock_get_s1_readdata;                   // clock_get:readdata -> mm_interconnect_0:clock_get_s1_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;       // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;           // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;             // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;              // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;          // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_btn_s1_writedata;                        // mm_interconnect_0:btn_s1_writedata -> btn:writedata
	wire   [1:0] mm_interconnect_0_btn_s1_address;                          // mm_interconnect_0:btn_s1_address -> btn:address
	wire         mm_interconnect_0_btn_s1_chipselect;                       // mm_interconnect_0:btn_s1_chipselect -> btn:chipselect
	wire         mm_interconnect_0_btn_s1_write;                            // mm_interconnect_0:btn_s1_write -> btn:write_n
	wire  [31:0] mm_interconnect_0_btn_s1_readdata;                         // btn:readdata -> mm_interconnect_0:btn_s1_readdata
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_writedata;     // mm_interconnect_0:lcd_16207_0_control_slave_writedata -> lcd_16207_0:writedata
	wire   [1:0] mm_interconnect_0_lcd_16207_0_control_slave_address;       // mm_interconnect_0:lcd_16207_0_control_slave_address -> lcd_16207_0:address
	wire         mm_interconnect_0_lcd_16207_0_control_slave_write;         // mm_interconnect_0:lcd_16207_0_control_slave_write -> lcd_16207_0:write
	wire         mm_interconnect_0_lcd_16207_0_control_slave_read;          // mm_interconnect_0:lcd_16207_0_control_slave_read -> lcd_16207_0:read
	wire   [7:0] mm_interconnect_0_lcd_16207_0_control_slave_readdata;      // lcd_16207_0:readdata -> mm_interconnect_0:lcd_16207_0_control_slave_readdata
	wire         mm_interconnect_0_lcd_16207_0_control_slave_begintransfer; // mm_interconnect_0:lcd_16207_0_control_slave_begintransfer -> lcd_16207_0:begintransfer
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire   [1:0] mm_interconnect_0_switch_s1_address;                       // mm_interconnect_0:switch_s1_address -> switch:address
	wire  [31:0] mm_interconnect_0_switch_s1_readdata;                      // switch:readdata -> mm_interconnect_0:switch_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire         mm_interconnect_0_sram_s1_waitrequest;                     // sram:za_waitrequest -> mm_interconnect_0:sram_s1_waitrequest
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                       // mm_interconnect_0:sram_s1_writedata -> sram:az_data
	wire  [23:0] mm_interconnect_0_sram_s1_address;                         // mm_interconnect_0:sram_s1_address -> sram:az_addr
	wire         mm_interconnect_0_sram_s1_chipselect;                      // mm_interconnect_0:sram_s1_chipselect -> sram:az_cs
	wire         mm_interconnect_0_sram_s1_write;                           // mm_interconnect_0:sram_s1_write -> sram:az_wr_n
	wire         mm_interconnect_0_sram_s1_read;                            // mm_interconnect_0:sram_s1_read -> sram:az_rd_n
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                        // sram:za_data -> mm_interconnect_0:sram_s1_readdata
	wire         mm_interconnect_0_sram_s1_readdatavalid;                   // sram:za_valid -> mm_interconnect_0:sram_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                      // mm_interconnect_0:sram_s1_byteenable -> sram:az_be_n
	wire         irq_mapper_receiver0_irq;                                  // btn:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // timer_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [btn:reset_n, clock_get:reset_n, clock_set:reset_n, cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, lcd_16207_0:reset_n, ledg:reset_n, ledr:reset_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sram:reset_n, switch:reset_n, sysid:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         clocks_sys_clk_reset_reset;                                // clocks:sys_reset_n -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> clocks:reset

	CPU_Final_Project_cpu cpu (
		.clk                                   (clocks_sys_clk_clk),                                  //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                    //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	CPU_Final_Project_sram sram (
		.clk            (clocks_sys_clk_clk),                      //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),         // reset.reset_n
		.az_addr        (mm_interconnect_0_sram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sram_wire_addr),                          //  wire.export
		.zs_ba          (sram_wire_ba),                            //      .export
		.zs_cas_n       (sram_wire_cas_n),                         //      .export
		.zs_cke         (sram_wire_cke),                           //      .export
		.zs_cs_n        (sram_wire_cs_n),                          //      .export
		.zs_dq          (sram_wire_dq),                            //      .export
		.zs_dqm         (sram_wire_dqm),                           //      .export
		.zs_ras_n       (sram_wire_ras_n),                         //      .export
		.zs_we_n        (sram_wire_we_n)                           //      .export
	);

	CPU_Final_Project_ledg ledg (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_external_connection_export)       // external_connection.export
	);

	CPU_Final_Project_ledr ledr (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)       // external_connection.export
	);

	CPU_Final_Project_switch switch (
		.clk      (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_s1_readdata), //                    .readdata
		.in_port  (switch_external_connection_export)     // external_connection.export
	);

	CPU_Final_Project_btn btn (
		.clk        (clocks_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_btn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_btn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_btn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_btn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_btn_s1_readdata),   //                    .readdata
		.in_port    (btn_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver0_irq)             //                 irq.irq
	);

	CPU_Final_Project_sysid sysid (
		.clock    (clocks_sys_clk_clk),                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	CPU_Final_Project_clocks clocks (
		.CLOCK_50    (clk_clk),                            //       clk_in_primary.clk
		.reset       (rst_controller_001_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (clocks_sys_clk_clk),                 //              sys_clk.clk
		.sys_reset_n (clocks_sys_clk_reset_reset),         //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clk_clk)                       //            sdram_clk.clk
	);

	CPU_Final_Project_lcd_16207_0 lcd_16207_0 (
		.reset_n       (~rst_controller_reset_out_reset),                           //         reset.reset_n
		.clk           (clocks_sys_clk_clk),                                        //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_16207_0_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_16207_0_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_16207_0_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_16207_0_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_16207_0_control_slave_address),       //              .address
		.LCD_RS        (lcd_16207_RS),                                              //      external.export
		.LCD_RW        (lcd_16207_RW),                                              //              .export
		.LCD_data      (lcd_16207_data),                                            //              .export
		.LCD_E         (lcd_16207_E)                                                //              .export
	);

	CPU_Final_Project_jtag_uart jtag_uart (
		.clk            (clocks_sys_clk_clk),                                        //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	CPU_Final_Project_clock_set clock_set (
		.clk        (clocks_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_clock_set_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_clock_set_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_clock_set_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_clock_set_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_clock_set_s1_readdata),   //                    .readdata
		.out_port   (clock_set_ext_export)                       // external_connection.export
	);

	CPU_Final_Project_clock_get clock_get (
		.clk      (clocks_sys_clk_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_clock_get_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_clock_get_s1_readdata), //                    .readdata
		.in_port  (clock_get_ext_export)                     // external_connection.export
	);

	CPU_Final_Project_timer_0 timer_0 (
		.clk        (clocks_sys_clk_clk),                      //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	CPU_Final_Project_mm_interconnect_0 mm_interconnect_0 (
		.clocks_sys_clk_clk                      (clocks_sys_clk_clk),                                        //                    clocks_sys_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                   cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                  .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                  .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                  .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                  .readdata
		.cpu_data_master_readdatavalid           (cpu_data_master_readdatavalid),                             //                                  .readdatavalid
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                  .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                  .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                  .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                  .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                  .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                  .readdata
		.cpu_instruction_master_readdatavalid    (cpu_instruction_master_readdatavalid),                      //                                  .readdatavalid
		.btn_s1_address                          (mm_interconnect_0_btn_s1_address),                          //                            btn_s1.address
		.btn_s1_write                            (mm_interconnect_0_btn_s1_write),                            //                                  .write
		.btn_s1_readdata                         (mm_interconnect_0_btn_s1_readdata),                         //                                  .readdata
		.btn_s1_writedata                        (mm_interconnect_0_btn_s1_writedata),                        //                                  .writedata
		.btn_s1_chipselect                       (mm_interconnect_0_btn_s1_chipselect),                       //                                  .chipselect
		.clock_get_s1_address                    (mm_interconnect_0_clock_get_s1_address),                    //                      clock_get_s1.address
		.clock_get_s1_readdata                   (mm_interconnect_0_clock_get_s1_readdata),                   //                                  .readdata
		.clock_set_s1_address                    (mm_interconnect_0_clock_set_s1_address),                    //                      clock_set_s1.address
		.clock_set_s1_write                      (mm_interconnect_0_clock_set_s1_write),                      //                                  .write
		.clock_set_s1_readdata                   (mm_interconnect_0_clock_set_s1_readdata),                   //                                  .readdata
		.clock_set_s1_writedata                  (mm_interconnect_0_clock_set_s1_writedata),                  //                                  .writedata
		.clock_set_s1_chipselect                 (mm_interconnect_0_clock_set_s1_chipselect),                 //                                  .chipselect
		.cpu_jtag_debug_module_address           (mm_interconnect_0_cpu_jtag_debug_module_address),           //             cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write             (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                  .write
		.cpu_jtag_debug_module_read              (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                  .read
		.cpu_jtag_debug_module_readdata          (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                  .readdata
		.cpu_jtag_debug_module_writedata         (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                  .writedata
		.cpu_jtag_debug_module_byteenable        (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                  .byteenable
		.cpu_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                  .waitrequest
		.cpu_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                  .debugaccess
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.lcd_16207_0_control_slave_address       (mm_interconnect_0_lcd_16207_0_control_slave_address),       //         lcd_16207_0_control_slave.address
		.lcd_16207_0_control_slave_write         (mm_interconnect_0_lcd_16207_0_control_slave_write),         //                                  .write
		.lcd_16207_0_control_slave_read          (mm_interconnect_0_lcd_16207_0_control_slave_read),          //                                  .read
		.lcd_16207_0_control_slave_readdata      (mm_interconnect_0_lcd_16207_0_control_slave_readdata),      //                                  .readdata
		.lcd_16207_0_control_slave_writedata     (mm_interconnect_0_lcd_16207_0_control_slave_writedata),     //                                  .writedata
		.lcd_16207_0_control_slave_begintransfer (mm_interconnect_0_lcd_16207_0_control_slave_begintransfer), //                                  .begintransfer
		.ledg_s1_address                         (mm_interconnect_0_ledg_s1_address),                         //                           ledg_s1.address
		.ledg_s1_write                           (mm_interconnect_0_ledg_s1_write),                           //                                  .write
		.ledg_s1_readdata                        (mm_interconnect_0_ledg_s1_readdata),                        //                                  .readdata
		.ledg_s1_writedata                       (mm_interconnect_0_ledg_s1_writedata),                       //                                  .writedata
		.ledg_s1_chipselect                      (mm_interconnect_0_ledg_s1_chipselect),                      //                                  .chipselect
		.ledr_s1_address                         (mm_interconnect_0_ledr_s1_address),                         //                           ledr_s1.address
		.ledr_s1_write                           (mm_interconnect_0_ledr_s1_write),                           //                                  .write
		.ledr_s1_readdata                        (mm_interconnect_0_ledr_s1_readdata),                        //                                  .readdata
		.ledr_s1_writedata                       (mm_interconnect_0_ledr_s1_writedata),                       //                                  .writedata
		.ledr_s1_chipselect                      (mm_interconnect_0_ledr_s1_chipselect),                      //                                  .chipselect
		.sram_s1_address                         (mm_interconnect_0_sram_s1_address),                         //                           sram_s1.address
		.sram_s1_write                           (mm_interconnect_0_sram_s1_write),                           //                                  .write
		.sram_s1_read                            (mm_interconnect_0_sram_s1_read),                            //                                  .read
		.sram_s1_readdata                        (mm_interconnect_0_sram_s1_readdata),                        //                                  .readdata
		.sram_s1_writedata                       (mm_interconnect_0_sram_s1_writedata),                       //                                  .writedata
		.sram_s1_byteenable                      (mm_interconnect_0_sram_s1_byteenable),                      //                                  .byteenable
		.sram_s1_readdatavalid                   (mm_interconnect_0_sram_s1_readdatavalid),                   //                                  .readdatavalid
		.sram_s1_waitrequest                     (mm_interconnect_0_sram_s1_waitrequest),                     //                                  .waitrequest
		.sram_s1_chipselect                      (mm_interconnect_0_sram_s1_chipselect),                      //                                  .chipselect
		.switch_s1_address                       (mm_interconnect_0_switch_s1_address),                       //                         switch_s1.address
		.switch_s1_readdata                      (mm_interconnect_0_switch_s1_readdata),                      //                                  .readdata
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //               sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata),            //                                  .readdata
		.timer_0_s1_address                      (mm_interconnect_0_timer_0_s1_address),                      //                        timer_0_s1.address
		.timer_0_s1_write                        (mm_interconnect_0_timer_0_s1_write),                        //                                  .write
		.timer_0_s1_readdata                     (mm_interconnect_0_timer_0_s1_readdata),                     //                                  .readdata
		.timer_0_s1_writedata                    (mm_interconnect_0_timer_0_s1_writedata),                    //                                  .writedata
		.timer_0_s1_chipselect                   (mm_interconnect_0_timer_0_s1_chipselect)                    //                                  .chipselect
	);

	CPU_Final_Project_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clocks_sys_clk_reset_reset),        // reset_in0.reset
		.clk            (clocks_sys_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
